<!DOCTYPE VIPEC_CIRCUIT_FILE  ><FILE VERSION="3.1.3" CREATOR="ViPEC" >
 <CIRCUIT SIZE="1" NAME="PRACTICARF4" >
  <COMPONENT TYPE="CLIN" >
   <LOCATION X="208" Y="120" ROTATION="0" />
   <TEXTOFFSET X="0" Y="0" />
   <ATTRIBUTE Ze="63.857" />
   <ATTRIBUTE Zo="51.468" />
   <ATTRIBUTE E="77.5715" />
   <ATTRIBUTE F="1.4" />
  </COMPONENT>
  <COMPONENT TYPE="PORT" >
   <LOCATION X="152" Y="112" ROTATION="0" />
   <TEXTOFFSET X="-1" Y="-29" />
   <ATTRIBUTE Z="50" />
  </COMPONENT>
  <COMPONENT TYPE="PORT" >
   <LOCATION X="272" Y="112" ROTATION="180" />
   <TEXTOFFSET X="3" Y="-31" />
   <ATTRIBUTE Z="50" />
  </COMPONENT>
  <COMPONENT TYPE="PORT" >
   <LOCATION X="152" Y="128" ROTATION="0" />
   <TEXTOFFSET X="0" Y="0" />
   <ATTRIBUTE Z="50" />
  </COMPONENT>
  <COMPONENT TYPE="PORT" >
   <LOCATION X="272" Y="128" ROTATION="180" />
   <TEXTOFFSET X="0" Y="0" />
   <ATTRIBUTE Z="50" />
  </COMPONENT>
  <LINE>
   <START X="160" Y="112" />
   <STOP X="184" Y="112" />
  </LINE>
  <LINE>
   <START X="264" Y="112" />
   <STOP X="232" Y="112" />
  </LINE>
  <LINE>
   <START X="160" Y="128" />
   <STOP X="184" Y="128" />
  </LINE>
  <LINE>
   <START X="264" Y="128" />
   <STOP X="232" Y="128" />
  </LINE>
 </CIRCUIT>
 <DIMENSIONS>
  <DIM VALUE="DEG" NAME="Angle" />
  <DIM VALUE="nF" NAME="Capacitance" />
  <DIM VALUE="GHz" NAME="Frequency" />
  <DIM VALUE="uH" NAME="Inductance" />
  <DIM VALUE="um" NAME="Length" />
  <DIM VALUE="Ohm" NAME="Resistance" />
  <DIM VALUE="us" NAME="Time" />
 </DIMENSIONS>
 <SWEEP STOP="3" POINTS="200" LINEAR="1" START="0.01" />
 <GRAPHDEFINITIONS>
  <GRID TITLE="1-2" NAME="PORT 1" >
   <XAXIS STEPS="5" MIN="0.01" MAX="3" TRACKING="1" />
   <YAXIS STEPS="5" MIN="-50" MAX="0" />
   <OUTPUT MEASUREMENT="0" DATASOURCE="PRACTICARF4" FORMAT="2" FROM="1" TYPE="0" TO="1" DB="1" />
   <OUTPUT MEASUREMENT="0" DATASOURCE="PRACTICARF4" FORMAT="2" FROM="2" TYPE="0" TO="1" DB="1" />
   <OUTPUT MEASUREMENT="0" DATASOURCE="PRACTICARF4" FORMAT="2" FROM="3" TYPE="0" TO="1" DB="1" />
   <OUTPUT MEASUREMENT="0" DATASOURCE="PRACTICARF4" FORMAT="2" FROM="4" TYPE="0" TO="1" DB="1" />
  </GRID>
  <GRID TITLE="" NAME="PORT 2" >
   <XAXIS STEPS="5" MIN="0.01" MAX="3" TRACKING="1" />
   <YAXIS STEPS="5" MIN="-50" MAX="0" />
   <OUTPUT MEASUREMENT="0" DATASOURCE="PRACTICARF4" FORMAT="2" FROM="2" TYPE="0" TO="2" DB="1" />
   <OUTPUT MEASUREMENT="0" DATASOURCE="PRACTICARF4" FORMAT="2" FROM="1" TYPE="0" TO="2" DB="1" />
   <OUTPUT MEASUREMENT="0" DATASOURCE="PRACTICARF4" FORMAT="2" FROM="3" TYPE="0" TO="2" DB="1" />
   <OUTPUT MEASUREMENT="0" DATASOURCE="PRACTICARF4" FORMAT="2" FROM="4" TYPE="0" TO="2" DB="1" />
  </GRID>
  <GRID TITLE="" NAME="PORT 3" >
   <XAXIS STEPS="5" MIN="0.01" MAX="3" TRACKING="1" />
   <YAXIS STEPS="5" MIN="-50" MAX="0" />
   <OUTPUT MEASUREMENT="0" DATASOURCE="PRACTICARF4" FORMAT="2" FROM="3" TYPE="0" TO="3" DB="1" />
   <OUTPUT MEASUREMENT="0" DATASOURCE="PRACTICARF4" FORMAT="2" FROM="1" TYPE="0" TO="3" DB="1" />
   <OUTPUT MEASUREMENT="0" DATASOURCE="PRACTICARF4" FORMAT="2" FROM="2" TYPE="0" TO="3" DB="1" />
   <OUTPUT MEASUREMENT="0" DATASOURCE="PRACTICARF4" FORMAT="2" FROM="4" TYPE="0" TO="3" DB="1" />
  </GRID>
  <GRID TITLE="" NAME="PORT 4" >
   <XAXIS STEPS="5" MIN="0.01" MAX="3" TRACKING="1" />
   <YAXIS STEPS="5" MIN="-50" MAX="0" />
   <OUTPUT MEASUREMENT="0" DATASOURCE="PRACTICARF4" FORMAT="2" FROM="4" TYPE="0" TO="4" DB="1" />
   <OUTPUT MEASUREMENT="0" DATASOURCE="PRACTICARF4" FORMAT="2" FROM="1" TYPE="0" TO="4" DB="1" />
   <OUTPUT MEASUREMENT="0" DATASOURCE="PRACTICARF4" FORMAT="2" FROM="2" TYPE="0" TO="4" DB="1" />
   <OUTPUT MEASUREMENT="0" DATASOURCE="PRACTICARF4" FORMAT="2" FROM="3" TYPE="0" TO="4" DB="1" />
  </GRID>
 </GRAPHDEFINITIONS>
 <SUBSTRATES/>
 <FILEBLOCKS/>
</FILE>
